Inverting OpAmp
* Inverting Op Amp
.lib eval.lib
.lib TL061.lib

*Vin 1 0 SIN(0 .1V 340Hz)
Vin 1 0 AC 1

Vcc 100 0 DC 9V

*RT1 2 0 10k

R1 3 4 2.7k
R2 3 5 10k

R3 100 9 100k
R4 9 0 100k
RT 9 2 10M

RL 6 0 100k

C1 4 0 10uF
C2 3 5 47pF
C3 5 6 1uF
C4 1 2 1uF
C5 9 0 1uF

X1 2 3 100 0 5 UA741

.TRAN 10nS .006S 0 5uS
.AC DEC 100 1HZ 5KHZ

.PROBE
.END

